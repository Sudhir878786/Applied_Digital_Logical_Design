`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    04:33:02 01/20/2020 
// Design Name: 
// Module Name:    addrev 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module addrev(
    input [3:0] a,
    input [3:0] b,
    output [3:0] c
    );

assign sum=a+b;

endmodule
